
// mem
`define ROM_ADDR_BASE		32'h0000_0000
`define ROM_SIZE		32'h0004_0000	// 128KB	
`define EF_BASE 		32'h1000_0000
`define EF_SIZE 		32'h1004_0000	// 256KB
`define SYSRAM_ADDR_BASE	32'h2000_0000
`define SYSRAM_SIZE		32'h0001_8000	// 64KB 
`define DATARAM_ADDR_BASE	32'h2002_0000
`define DATARAM_SIZE		32'h0000_2000	// 8KB

// io
`define REG_SIZE		32'h0000_0100	// 256B
`define BLE_REG_SIZE		32'h0002_0000	// 8k use 16k
`define SCU_ADDR_BASE		32'h4000_0000
`define CKGEN_ADDR_BASE		32'h4000_0100
`define GPIO_ADDR_BASE		32'h4000_0200
`define WDT_ADDR_BASE		32'h4000_0300
`define PWM0_ADDR_BASE		32'h4000_0400
`define PWM1_ADDR_BASE		32'h4000_0500
`define WKTM0_ADDR_BASE		32'h4000_0600
`define WKTM1_ADDR_BASE		32'h4000_0700

`define RTC_ADDR_BASE		32'h4000_0800
`define I2S_ADDR_BASE		32'h4000_0900
`define DMIC_ADDR_BASE		32'h4000_0a00
`define SPI0_ADDR_BASE		32'h4000_0b00
`define SPI1_ADDR_BASE		32'h4000_0c00
`define SPI2_ADDR_BASE		32'h4000_0d00
`define UART0_ADDR_BASE		32'h4000_0e00
`define UART1_ADDR_BASE		32'h4000_0f00
	
`define UART2_ADDR_BASE		32'h4000_1000
`define I2C0_ADDR_BASE		32'h4000_1100
`define I2C1_ADDR_BASE		32'h4000_1200
`define DMU_ADDR_BASE		32'h4000_1300

`define EF_ADDR_BASE		32'h4000_2000
`define OTP_ADDR_BASE		32'h4000_2100
`define HS_ADDR_BASE		32'h4000_2200
`define PMU_ADDR_BASE		32'h4000_2300
`define AES_ADDR_BASE		32'h4000_2400
`define CCU_ADDR_BASE		32'h4000_2500

`define BLE_ADDR_BASE		32'h4000_4000

// EF
`define EF_INTERRUPT_REG   `EF_ADDR_BASE + 32'h0000_0000
`define EF_CONFIG_REG      `EF_ADDR_BASE + 32'h0000_0004
`define EF_ACCESS_REG      `EF_ADDR_BASE + 32'h0000_0008
`define EF_WR_DATA0_REG    `EF_ADDR_BASE + 32'h0000_000c
`define EF_WR_DATA1_REG    `EF_ADDR_BASE + 32'h0000_0010
`define EF_WR_DATA2_REG    `EF_ADDR_BASE + 32'h0000_0014
`define EF_WR_DATA3_REG    `EF_ADDR_BASE + 32'h0000_0018
`define EF_FLASHMODE_REG   `EF_ADDR_BASE + 32'h0000_001c
`define EF_RD_DATA0_REG    `EF_ADDR_BASE + 32'h0000_0020
`define EF_RD_DATA1_REG    `EF_ADDR_BASE + 32'h0000_0024
`define EF_REDUN_DATA_REG  `EF_ADDR_BASE + 32'h0000_0028

`define EF_TIMING0_REG     `EF_ADDR_BASE + 32'h0000_0044
`define EF_TIMING1_REG     `EF_ADDR_BASE + 32'h0000_0048
`define EF_TIMING2_REG     `EF_ADDR_BASE + 32'h0000_004c
`define EF_TIMING3_REG     `EF_ADDR_BASE + 32'h0000_0050
`define EF_TIMING4_REG     `EF_ADDR_BASE + 32'h0000_0054
`define EF_TIMING5_REG     `EF_ADDR_BASE + 32'h0000_0058
`define EF_TIMING6_REG     `EF_ADDR_BASE + 32'h0000_005c

`define EF_DMA_CTRL_REG	   `EF_ADDR_BASE + 32'h0000_0060
`define EF_DMA_WADDR_REG   `EF_ADDR_BASE + 32'h0000_0064
`define EF_DMA_RADDR_REG   `EF_ADDR_BASE + 32'h0000_0068

// SCU
`define SCU_INTRCTRL_REG	`SCU_ADDR_BASE + 32'h0000_0000
`define SCU_PLLLOCK_REG		`SCU_ADDR_BASE + 32'h0000_0004
`define SCU_PLLRST_REG		`SCU_ADDR_BASE + 32'h0000_0008
`define SCU_PLLCFG_REG		`SCU_ADDR_BASE + 32'h0000_000c
`define SCU_CLKCFG0_REG		`SCU_ADDR_BASE + 32'h0000_0010
`define SCU_CLKCFG1_REG		`SCU_ADDR_BASE + 32'h0000_0014
`define SCU_CHIPID_REG		`SCU_ADDR_BASE + 32'h0000_001c
`define SCU_ISOCTRL_REG		`SCU_ADDR_BASE + 32'h0000_0020
`define SCU_PSOCTRL_REG		`SCU_ADDR_BASE + 32'h0000_0024
`define SCU_RETCTRL_REG		`SCU_ADDR_BASE + 32'h0000_0028
`define SCU_EXTAUX_REG		`SCU_ADDR_BASE + 32'h0000_002c
`define SCU_HSCLK_REG		`SCU_ADDR_BASE + 32'h0000_0030
`define SCU_ICACHE_REG		`SCU_ADDR_BASE + 32'h0000_0034
`define SCU_CLK32K_CAL_REG	`SCU_ADDR_BASE + 32'h0000_0038
`define SCU_INTRMASK_REG	`SCU_ADDR_BASE + 32'h0000_003c
`define SCU_INTRINFO_REG	`SCU_ADDR_BASE + 32'h0000_0040	

// CKGEN
`define CKGEN_CFG1_REG		`CKGEN_ADDR_BASE + 32'h0000_0004
`define CKGEN_CFG2_REG		`CKGEN_ADDR_BASE + 32'h0000_0008
`define CKGEN_CFG3_REG		`CKGEN_ADDR_BASE + 32'h0000_000c
`define CKGEN_CFG4_REG		`CKGEN_ADDR_BASE + 32'h0000_0010
`define CKGEN_CLKEN_REG		`CKGEN_ADDR_BASE + 32'h0000_0014
`define CKGEN_SWRST_REG   	`CKGEN_ADDR_BASE + 32'h0000_0018
`define CKGEN_BLECLKSEL_REG 	`CKGEN_ADDR_BASE + 32'h0000_001c

// GPIO
`define GPIO_PAD_OUT_REG	`GPIO_ADDR_BASE + 32'h0000_0000
`define GPIO_PAD_IN_REG		`GPIO_ADDR_BASE + 32'h0000_0004
`define GPIO_PAD_OE_REG		`GPIO_ADDR_BASE + 32'h0000_0008
`define GPIO_INTR_PRIO_REG	`GPIO_ADDR_BASE + 32'h0000_000c
`define GPIO_INTR_EN_REG	`GPIO_ADDR_BASE + 32'h0000_0010
`define GPIO_INTR_STAT_REG	`GPIO_ADDR_BASE + 32'h0000_0014
`define GPIO_INTR_TRIG_REG	`GPIO_ADDR_BASE + 32'h0000_0018
`define GPIO_AUX_REG		`GPIO_ADDR_BASE + 32'h0000_001c
`define GPIO_INTR_TYPE_REG	`GPIO_ADDR_BASE + 32'h0000_0020
`define GPIO_PAD_PULLUP_REG	`GPIO_ADDR_BASE + 32'h0000_0024
`define GPIO_AUX_PORT_MODE_REG	`GPIO_ADDR_BASE + 32'h0000_0028

`define GPIO1_PAD_OUT_REG       `GPIO_ADDR_BASE + 32'h0000_002c
`define GPIO1_PAD_IN_REG        `GPIO_ADDR_BASE + 32'h0000_0030
`define GPIO1_PAD_OE_REG        `GPIO_ADDR_BASE + 32'h0000_0034
`define GPIO1_INTR_PRIO_REG     `GPIO_ADDR_BASE + 32'h0000_0038
`define GPIO1_INTR_EN_REG       `GPIO_ADDR_BASE + 32'h0000_003c
`define GPIO1_INTR_STAT_REG     `GPIO_ADDR_BASE + 32'h0000_0040
`define GPIO1_INTR_TRIG_REG     `GPIO_ADDR_BASE + 32'h0000_0044
`define GPIO1_AUX_REG           `GPIO_ADDR_BASE + 32'h0000_0048
`define GPIO1_INTR_TYPE_REG     `GPIO_ADDR_BASE + 32'h0000_004c
`define GPIO1_PAD_PULLUP_REG    `GPIO_ADDR_BASE + 32'h0000_0050
`define GPIO1_AUX_PORT_MODE_REG `GPIO_ADDR_BASE + 32'h0000_0054

// SPI
`define SPI0_INTR_REG		`SPI0_ADDR_BASE + 32'h0000_0000
`define SPI0_CTRL_REG		`SPI0_ADDR_BASE + 32'h0000_0004
`define SPI0_DMA_CTRL_REG	`SPI0_ADDR_BASE + 32'h0000_0008
`define SPI0_DMA_WR_REG		`SPI0_ADDR_BASE + 32'h0000_000c
`define SPI0_DMA_RD_REG		`SPI0_ADDR_BASE + 32'h0000_0010

`define SPI1_INTR_REG           `SPI1_ADDR_BASE + 32'h0000_0000
`define SPI1_CTRL_REG           `SPI1_ADDR_BASE + 32'h0000_0004
`define SPI1_DMA_CTRL_REG       `SPI1_ADDR_BASE + 32'h0000_0008
`define SPI1_DMA_WR_REG         `SPI1_ADDR_BASE + 32'h0000_000c
`define SPI1_DMA_RD_REG         `SPI1_ADDR_BASE + 32'h0000_0010

`define SPI1_INTR_REG           `SPI1_ADDR_BASE + 32'h0000_0000
`define SPI1_CTRL_REG           `SPI1_ADDR_BASE + 32'h0000_0004
`define SPI1_DMA_CTRL_REG       `SPI1_ADDR_BASE + 32'h0000_0008
`define SPI1_DMA_WR_REG         `SPI1_ADDR_BASE + 32'h0000_000c
`define SPI1_DMA_RD_REG         `SPI1_ADDR_BASE + 32'h0000_0010

// WDT
`define WDT_TIMER0_REG		`WDT_ADDR_BASE + 32'h0000_0000
`define WDT_TIMER1_REG		`WDT_ADDR_BASE + 32'h0000_0004
`define WDT_TIMER2_REG		`WDT_ADDR_BASE + 32'h0000_0008
`define WDT_TIMER3_REG		`WDT_ADDR_BASE + 32'h0000_000c

// RTC
`define RTC_SEC_REG		`RTC_ADDR_BASE + 32'h0000_0000
`define RTC_MIN_REG		`RTC_ADDR_BASE + 32'h0000_0004
`define RTC_HRS_REG		`RTC_ADDR_BASE + 32'h0000_0008
`define RTC_DOW_REG		`RTC_ADDR_BASE + 32'h0000_000c
`define RTC_DAY_REG		`RTC_ADDR_BASE + 32'h0000_0010
`define RTC_MON_REG		`RTC_ADDR_BASE + 32'h0000_0014
`define RTC_YRS_REG		`RTC_ADDR_BASE + 32'h0000_0018

`define RTC_ALM_SEC_REG		`RTC_ADDR_BASE + 32'h0000_001c
`define RTC_ALM_MIN_REG		`RTC_ADDR_BASE + 32'h0000_0020
`define RTC_ALM_HRS_REG		`RTC_ADDR_BASE + 32'h0000_0024
`define RTC_ALM_DOM_REG		`RTC_ADDR_BASE + 32'h0000_0028
`define RTC_ALM_MON_REG		`RTC_ADDR_BASE + 32'h0000_002c

`define RTC_ALM2_SEC_REG        `RTC_ADDR_BASE + 32'h0000_0030
`define RTC_ALM2_MIN_REG        `RTC_ADDR_BASE + 32'h0000_0034
`define RTC_ALM2_HRS_REG        `RTC_ADDR_BASE + 32'h0000_0038
`define RTC_ALM2_DOM_REG        `RTC_ADDR_BASE + 32'h0000_003c
`define RTC_ALM2_MON_REG        `RTC_ADDR_BASE + 32'h0000_0040

`define RTC_CTRLA_REG		`RTC_ADDR_BASE + 32'h0000_0044
`define RTC_CTRLB_REG		`RTC_ADDR_BASE + 32'h0000_0048
`define RTC_CTRLC_REG		`RTC_ADDR_BASE + 32'h0000_0050

// CCU
`define CCU_INTR_REG		`CCU_ADDR_BASE + 32'h0000_0000
`define CCU_DELTA_CNT_REG	`CCU_ADDR_BASE + 32'h0000_0004
`define CCU_FDELTA_CNT_REG	`CCU_ADDR_BASE + 32'h0000_0008

// UART
`define UART0_UnBAUD_REG	`UART0_ADDR_BASE + 32'h0000_0018
`define UART0_UnPSR_REG		`UART0_ADDR_BASE + 32'h0000_001c
`define UART0_UnOVR_REG		`UART0_ADDR_BASE + 32'h0000_0020

`define UART1_UnBAUD_REG        `UART1_ADDR_BASE + 32'h0000_0018
`define UART1_UnPSR_REG         `UART1_ADDR_BASE + 32'h0000_001c
`define UART1_UnOVR_REG         `UART1_ADDR_BASE + 32'h0000_0020

`define UART2_UnBAUD_REG        `UART2_ADDR_BASE + 32'h0000_0018
`define UART2_UnPSR_REG         `UART2_ADDR_BASE + 32'h0000_001c
`define UART2_UnOVR_REG         `UART2_ADDR_BASE + 32'h0000_0020

// HS
`define HS_CONFIG_REG		`HS_ADDR_BASE + 32'h0000_0000
`define HS_STS_REG		`HS_ADDR_BASE + 32'h0000_0004
`define HS_DR_PDN_REG		`HS_ADDR_BASE + 32'h0000_0008
`define HS_DR0_PUP_REG		`HS_ADDR_BASE + 32'h0000_000c
`define HS_DR0_PUP1_REG		`HS_ADDR_BASE + 32'h0000_0010
`define HS_DR0_INTR_REG		`HS_ADDR_BASE + 32'h0000_0014
`define HS_DR1_PUP_REG          `HS_ADDR_BASE + 32'h0000_0018
`define HS_DR1_PUP1_REG         `HS_ADDR_BASE + 32'h0000_001c
`define HS_DR1_INTR_REG		`HS_ADDR_BASE + 32'h0000_0020
`define HS_DR2_PUP_REG          `HS_ADDR_BASE + 32'h0000_0024
`define HS_DR2_PUP1_REG         `HS_ADDR_BASE + 32'h0000_0028
`define HS_DR2_INTR_REG		`HS_ADDR_BASE + 32'h0000_002c
`define HS_SCRATCH_BASE_REG	`HS_ADDR_BASE + 32'h0000_0030

// INTERRUPT
`define EF_INTR 		`CHIP_CORE0.interrupt_o[31]
`define SPI0_EXT_INTR		`CHIP_CORE0.interrupt_o[30]
`define I2C0_EXT_INTR		`CHIP_CORE0.interrupt_o[29]
`define AES_INTR		`CHIP_CORE0.interrupt_o[28]
`define CCU_INTR		`CHIP_CORE0.interrupt_o[27]
`define GPIO_INTR		`CHIP_CORE0.interrupt_o[26]
`define BLE_INTR		`CHIP_CORE0.interrupt_o[25]
`define DMIC_INTR		`CHIP_CORE0.interrupt_o[24]
`define I2S_IP_INTR		`CHIP_CORE0.interrupt_o[23]
`define I2S_TXDMA_INTR		`CHIP_CORE0.interrupt_o[22]
`define I2S_RXDMA_INTR		`CHIP_CORE0.interrupt_o[21]
`define I2C1_INTR		`CHIP_CORE0.interrupt_o[20]
`define I2C0_INTR		`CHIP_CORE0.interrupt_o[19]
`define UART2_IP_INTR		`CHIP_CORE0.interrupt_o[18]
`define UART2_TXDMA_INTR	`CHIP_CORE0.interrupt_o[17]
`define UART2_RXDMA_INTR	`CHIP_CORE0.interrupt_o[16]
`define UART1_IP_INTR   	`CHIP_CORE0.interrupt_o[15]
`define UART1_TXDMA_INTR        `CHIP_CORE0.interrupt_o[14]
`define UART1_RXDMA_INTR        `CHIP_CORE0.interrupt_o[13]
`define UART0_IP_INTR   	`CHIP_CORE0.interrupt_o[12]
`define UART0_TXDMA_INTR        `CHIP_CORE0.interrupt_o[11]
`define UART0_RXDMA_INTR        `CHIP_CORE0.interrupt_o[10]
`define	SPI2_M_INTR		`CHIP_CORE0.interrupt_o[9]
`define SPI1_M_INTR		`CHIP_CORE0.interrupt_o[8]
`define SPI0_M_INTR		`CHIP_CORE0.interrupt_o[7]
`define WKT1_INTR		`CHIP_CORE0.interrupt_o[6]
`define WKT0_INTR		`CHIP_CORE0.interrupt_o[5]
`define PWM1_INTR		`CHIP_CORE0.interrupt_o[4]
`define PWM0_INTR		`CHIP_CORE0.interrupt_o[3]
`define RTC_INTR		`CHIP_CORE0.interrupt_o[2]
`define WDT_INTR		`CHIP_CORE0.interrupt_o[1]
`define SCU_INTR		`CHIP_CORE0.interrupt_o[0]



